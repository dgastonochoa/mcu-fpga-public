`ifndef TEST_MCU_SVH
`define TEST_MCU_SVH

`define MCU_GET_M(mcu) mcu.cm
`define MCU_GET_C(mcu) mcu.c

`endif // TEST_MCU_SVH