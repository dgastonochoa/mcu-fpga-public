`ifndef RISCV_SINGLE_ALL_INSTR_MEM_MAP_SVH
`define RISCV_SINGLE_ALL_INSTR_MEM_MAP_SVH
/**
 * This file is to be used by the @see{mem.sv} module if
 * CONFIG_ENABLE_MEM_DEFAULT_VALS is enabled.
 */

`define INIT_MEM_F(mem_reg)         \
    mem_reg[0] = 32'h6c000113;      \
    mem_reg[1] = 32'h02500293;      \
    mem_reg[2] = 32'h00328313;      \
    mem_reg[3] = 32'h00512023;      \
    mem_reg[4] = 32'h00612223;      \
    mem_reg[5] = 32'h004001ef;      \
    mem_reg[6] = 32'h00312423;      \
    mem_reg[7] = 32'habcde2b7;      \
    mem_reg[8] = 32'h00f12337;      \
    mem_reg[9] = 32'h00c35313;      \
    mem_reg[10] = 32'h0062e2b3;     \
    mem_reg[11] = 32'h00512623;     \
    mem_reg[12] = 32'h00000293;     \
    mem_reg[13] = 32'h00c14283;     \
    mem_reg[14] = 32'h00512823;     \
    mem_reg[15] = 32'h00000293;     \
    mem_reg[16] = 32'h00d14283;     \
    mem_reg[17] = 32'h00512a23;     \
    mem_reg[18] = 32'h00000293;     \
    mem_reg[19] = 32'h00e14283;     \
    mem_reg[20] = 32'h00512c23;     \
    mem_reg[21] = 32'h00000293;     \
    mem_reg[22] = 32'h00f14283;     \
    mem_reg[23] = 32'h00512e23;     \
    mem_reg[24] = 32'h00000293;     \
    mem_reg[25] = 32'h00c15283;     \
    mem_reg[26] = 32'h02512023;     \
    mem_reg[27] = 32'h00000293;     \
    mem_reg[28] = 32'h00e15283;     \
    mem_reg[29] = 32'h02512223;     \
    mem_reg[30] = 32'h00000293;     \
    mem_reg[31] = 32'h00c12283;     \
    mem_reg[32] = 32'h02512423;     \
    mem_reg[33] = 32'h02511623;     \
    mem_reg[34] = 32'h02510823;     \
    mem_reg[35] = 32'h00000293;     \
    mem_reg[36] = 32'h00c10283;     \
    mem_reg[37] = 32'h02512a23;     \
    mem_reg[38] = 32'h00000293;     \
    mem_reg[39] = 32'h00d10283;     \
    mem_reg[40] = 32'h02512c23;     \
    mem_reg[41] = 32'h00000293;     \
    mem_reg[42] = 32'h00e10283;     \
    mem_reg[43] = 32'h02512e23;     \
    mem_reg[44] = 32'h00000293;     \
    mem_reg[45] = 32'h00f10283;     \
    mem_reg[46] = 32'h04512023;     \
    mem_reg[47] = 32'h00000293;     \
    mem_reg[48] = 32'h00c11283;     \
    mem_reg[49] = 32'h04512223;     \
    mem_reg[50] = 32'h00000293;     \
    mem_reg[51] = 32'h7ffff2b7;     \
    mem_reg[52] = 32'h04512423;     \
    mem_reg[53] = 32'h00000293;     \
    mem_reg[54] = 32'h04a11283;     \
    mem_reg[55] = 32'h00c12283;     \
    mem_reg[56] = 32'h00829313;     \
    mem_reg[57] = 32'h04612623;     \
    mem_reg[58] = 32'h00929313;     \
    mem_reg[59] = 32'h04612823;     \
    mem_reg[60] = 32'h00029313;     \
    mem_reg[61] = 32'h04612a23;     \
    mem_reg[62] = 32'h01f29313;     \
    mem_reg[63] = 32'h04612c23;     \
    mem_reg[64] = 32'h00700313;     \
    mem_reg[65] = 32'h00632393;     \
    mem_reg[66] = 32'h04712e23;     \
    mem_reg[67] = 32'h00832393;     \
    mem_reg[68] = 32'h06712023;     \
    mem_reg[69] = 32'hffd32393;     \
    mem_reg[70] = 32'h06712223;     \
    mem_reg[71] = 32'h00032393;     \
    mem_reg[72] = 32'h06712423;     \
    mem_reg[73] = 32'h00732393;     \
    mem_reg[74] = 32'h06712623;     \
    mem_reg[75] = 32'h00000313;     \
    mem_reg[76] = 32'h00632393;     \
    mem_reg[77] = 32'h06712823;     \
    mem_reg[78] = 32'hffd32393;     \
    mem_reg[79] = 32'h06712a23;     \
    mem_reg[80] = 32'h00032393;     \
    mem_reg[81] = 32'h06712c23;     \
    mem_reg[82] = 32'hff900313;     \
    mem_reg[83] = 32'hff832393;     \
    mem_reg[84] = 32'h06712e23;     \
    mem_reg[85] = 32'hff932393;     \
    mem_reg[86] = 32'h08712023;     \
    mem_reg[87] = 32'hffa32393;     \
    mem_reg[88] = 32'h08712223;     \
    mem_reg[89] = 32'h00032393;     \
    mem_reg[90] = 32'h08712423;     \
    mem_reg[91] = 32'h00832393;     \
    mem_reg[92] = 32'h08712623;     \
    mem_reg[93] = 32'h00700313;     \
    mem_reg[94] = 32'h00633393;     \
    mem_reg[95] = 32'h08712823;     \
    mem_reg[96] = 32'h00833393;     \
    mem_reg[97] = 32'h08712a23;     \
    mem_reg[98] = 32'hffd33393;     \
    mem_reg[99] = 32'h08712c23;     \
    mem_reg[100] = 32'h00033393;        \
    mem_reg[101] = 32'h08712e23;        \
    mem_reg[102] = 32'h00733393;        \
    mem_reg[103] = 32'h0a712023;        \
    mem_reg[104] = 32'h00000313;        \
    mem_reg[105] = 32'h00633393;        \
    mem_reg[106] = 32'h0a712223;        \
    mem_reg[107] = 32'hffd33393;        \
    mem_reg[108] = 32'h0a712423;        \
    mem_reg[109] = 32'h00033393;        \
    mem_reg[110] = 32'h0a712623;        \
    mem_reg[111] = 32'hff900313;        \
    mem_reg[112] = 32'hff833393;        \
    mem_reg[113] = 32'h0a712823;        \
    mem_reg[114] = 32'hff933393;        \
    mem_reg[115] = 32'h0a712a23;        \
    mem_reg[116] = 32'hffa33393;        \
    mem_reg[117] = 32'h0a712c23;        \
    mem_reg[118] = 32'h00033393;        \
    mem_reg[119] = 32'h0a712e23;        \
    mem_reg[120] = 32'h00833393;        \
    mem_reg[121] = 32'h0c712023;        \
    mem_reg[122] = 32'h0aa00313;        \
    mem_reg[123] = 32'h05534393;        \
    mem_reg[124] = 32'h0c712223;        \
    mem_reg[125] = 32'h0ff3c393;        \
    mem_reg[126] = 32'h0c712423;        \
    mem_reg[127] = 32'hfffff337;        \
    mem_reg[128] = 32'h00435393;        \
    mem_reg[129] = 32'h0c712623;        \
    mem_reg[130] = 32'h00835393;        \
    mem_reg[131] = 32'h0c712823;        \
    mem_reg[132] = 32'hfffff337;        \
    mem_reg[133] = 32'h40435393;        \
    mem_reg[134] = 32'h0c712a23;        \
    mem_reg[135] = 32'h40835393;        \
    mem_reg[136] = 32'h0c712c23;        \
    mem_reg[137] = 32'h00000313;        \
    mem_reg[138] = 32'h0f036393;        \
    mem_reg[139] = 32'h0c712e23;        \
    mem_reg[140] = 32'h0ff36393;        \
    mem_reg[141] = 32'h0e712023;        \
    mem_reg[142] = 32'h0003e393;        \
    mem_reg[143] = 32'h0e712223;        \
    mem_reg[144] = 32'h7ff00313;        \
    mem_reg[145] = 32'h0ff37393;        \
    mem_reg[146] = 32'h0e712423;        \
    mem_reg[147] = 32'h00f37393;        \
    mem_reg[148] = 32'h0e712623;        \
    mem_reg[149] = 32'h00037393;        \
    mem_reg[150] = 32'h0e712823;        \
    mem_reg[151] = 32'h00001317;        \
    mem_reg[152] = 32'h00001397;        \
    mem_reg[153] = 32'h406383b3;        \
    mem_reg[154] = 32'h0e712a23;        \
    mem_reg[155] = 32'h00c12283;        \
    mem_reg[156] = 32'h00800413;        \
    mem_reg[157] = 32'h00829333;        \
    mem_reg[158] = 32'h0e612c23;        \
    mem_reg[159] = 32'h00900413;        \
    mem_reg[160] = 32'h00829333;        \
    mem_reg[161] = 32'h0e612e23;        \
    mem_reg[162] = 32'h00000413;        \
    mem_reg[163] = 32'h00829333;        \
    mem_reg[164] = 32'h10612023;        \
    mem_reg[165] = 32'h01f00413;        \
    mem_reg[166] = 32'h00829333;        \
    mem_reg[167] = 32'h10612223;        \
    mem_reg[168] = 32'h00700313;        \
    mem_reg[169] = 32'h00600413;        \
    mem_reg[170] = 32'h008323b3;        \
    mem_reg[171] = 32'h10712223;        \
    mem_reg[172] = 32'h00800413;        \
    mem_reg[173] = 32'h008323b3;        \
    mem_reg[174] = 32'h10712423;        \
    mem_reg[175] = 32'hffd00413;        \
    mem_reg[176] = 32'h008323b3;        \
    mem_reg[177] = 32'h10712623;        \
    mem_reg[178] = 32'h00000413;        \
    mem_reg[179] = 32'h008323b3;        \
    mem_reg[180] = 32'h10712823;        \
    mem_reg[181] = 32'h00700413;        \
    mem_reg[182] = 32'h008323b3;        \
    mem_reg[183] = 32'h10712a23;        \
    mem_reg[184] = 32'h00000313;        \
    mem_reg[185] = 32'h00600413;        \
    mem_reg[186] = 32'h008323b3;        \
    mem_reg[187] = 32'h10712c23;        \
    mem_reg[188] = 32'hffd00413;        \
    mem_reg[189] = 32'h008323b3;        \
    mem_reg[190] = 32'h10712e23;        \
    mem_reg[191] = 32'h00000413;        \
    mem_reg[192] = 32'h008323b3;        \
    mem_reg[193] = 32'h12712023;        \
    mem_reg[194] = 32'hff900313;        \
    mem_reg[195] = 32'hff800413;        \
    mem_reg[196] = 32'h008323b3;        \
    mem_reg[197] = 32'h12712223;        \
    mem_reg[198] = 32'hff900413;        \
    mem_reg[199] = 32'h008323b3;        \
    mem_reg[200] = 32'h12712423;        \
    mem_reg[201] = 32'hffa00413;        \
    mem_reg[202] = 32'h008323b3;        \
    mem_reg[203] = 32'h12712623;        \
    mem_reg[204] = 32'h00000413;        \
    mem_reg[205] = 32'h008323b3;        \
    mem_reg[206] = 32'h12712823;        \
    mem_reg[207] = 32'h00800413;        \
    mem_reg[208] = 32'h008323b3;        \
    mem_reg[209] = 32'h12712a23;        \
    mem_reg[210] = 32'h00700313;        \
    mem_reg[211] = 32'h00600413;        \
    mem_reg[212] = 32'h008333b3;        \
    mem_reg[213] = 32'h12712c23;        \
    mem_reg[214] = 32'h00800413;        \
    mem_reg[215] = 32'h008333b3;        \
    mem_reg[216] = 32'h12712e23;        \
    mem_reg[217] = 32'hffd00413;        \
    mem_reg[218] = 32'h008333b3;        \
    mem_reg[219] = 32'h14712023;        \
    mem_reg[220] = 32'h00000413;        \
    mem_reg[221] = 32'h008333b3;        \
    mem_reg[222] = 32'h14712223;        \
    mem_reg[223] = 32'h00700413;        \
    mem_reg[224] = 32'h008333b3;        \
    mem_reg[225] = 32'h14712423;        \
    mem_reg[226] = 32'h00000313;        \
    mem_reg[227] = 32'h00600413;        \
    mem_reg[228] = 32'h008333b3;        \
    mem_reg[229] = 32'h14712623;        \
    mem_reg[230] = 32'hffd00413;        \
    mem_reg[231] = 32'h008333b3;        \
    mem_reg[232] = 32'h14712823;        \
    mem_reg[233] = 32'h00000413;        \
    mem_reg[234] = 32'h008333b3;        \
    mem_reg[235] = 32'h14712a23;        \
    mem_reg[236] = 32'hff900313;        \
    mem_reg[237] = 32'hff800413;        \
    mem_reg[238] = 32'h008333b3;        \
    mem_reg[239] = 32'h14712c23;        \
    mem_reg[240] = 32'hff900413;        \
    mem_reg[241] = 32'h008333b3;        \
    mem_reg[242] = 32'h14712e23;        \
    mem_reg[243] = 32'hffa00413;        \
    mem_reg[244] = 32'h008333b3;        \
    mem_reg[245] = 32'h16712023;        \
    mem_reg[246] = 32'h00000413;        \
    mem_reg[247] = 32'h008333b3;        \
    mem_reg[248] = 32'h16712223;        \
    mem_reg[249] = 32'h00800413;        \
    mem_reg[250] = 32'h008333b3;        \
    mem_reg[251] = 32'h16712423;        \
    mem_reg[252] = 32'h0aa00313;        \
    mem_reg[253] = 32'h05500413;        \
    mem_reg[254] = 32'h008343b3;        \
    mem_reg[255] = 32'h16712623;        \
    mem_reg[256] = 32'h0ff00413;        \
    mem_reg[257] = 32'h0083c3b3;        \
    mem_reg[258] = 32'h16712823;        \
    mem_reg[259] = 32'hfffff337;        \
    mem_reg[260] = 32'h00400413;        \
    mem_reg[261] = 32'h008353b3;        \
    mem_reg[262] = 32'h16712a23;        \
    mem_reg[263] = 32'h00800413;        \
    mem_reg[264] = 32'h008353b3;        \
    mem_reg[265] = 32'h16712c23;        \
    mem_reg[266] = 32'hfffff337;        \
    mem_reg[267] = 32'h00400413;        \
    mem_reg[268] = 32'h408353b3;        \
    mem_reg[269] = 32'h16712e23;        \
    mem_reg[270] = 32'h00800413;        \
    mem_reg[271] = 32'h408353b3;        \
    mem_reg[272] = 32'h18712023;        \
    mem_reg[273] = 32'h00000313;        \
    mem_reg[274] = 32'h0f000413;        \
    mem_reg[275] = 32'h008363b3;        \
    mem_reg[276] = 32'h18712223;        \
    mem_reg[277] = 32'h0ff00413;        \
    mem_reg[278] = 32'h008363b3;        \
    mem_reg[279] = 32'h18712423;        \
    mem_reg[280] = 32'h00000413;        \
    mem_reg[281] = 32'h0083e3b3;        \
    mem_reg[282] = 32'h18712623;        \
    mem_reg[283] = 32'h7ff00313;        \
    mem_reg[284] = 32'h0ff00413;        \
    mem_reg[285] = 32'h008373b3;        \
    mem_reg[286] = 32'h18712823;        \
    mem_reg[287] = 32'h00f00413;        \
    mem_reg[288] = 32'h008373b3;        \
    mem_reg[289] = 32'h18712a23;        \
    mem_reg[290] = 32'h00000413;        \
    mem_reg[291] = 32'h008373b3;        \
    mem_reg[292] = 32'h18712c23;        \
    mem_reg[293] = 32'h01400313;        \
    mem_reg[294] = 32'h00030393;        \
    mem_reg[295] = 32'h18712e23;        \
    mem_reg[296] = 32'h00530393;        \
    mem_reg[297] = 32'h1a712023;        \
    mem_reg[298] = 32'hfec30393;        \
    mem_reg[299] = 32'h1a712223;        \
    mem_reg[300] = 32'hfe730393;        \
    mem_reg[301] = 32'h1a712423;        \
    mem_reg[302] = 32'h01400313;        \
    mem_reg[303] = 32'h00000413;        \
    mem_reg[304] = 32'h008303b3;        \
    mem_reg[305] = 32'h1a712623;        \
    mem_reg[306] = 32'h00500413;        \
    mem_reg[307] = 32'h008303b3;        \
    mem_reg[308] = 32'h1a712823;        \
    mem_reg[309] = 32'hfec00413;        \
    mem_reg[310] = 32'h008303b3;        \
    mem_reg[311] = 32'h1a712a23;        \
    mem_reg[312] = 32'hfe700413;        \
    mem_reg[313] = 32'h008303b3;        \
    mem_reg[314] = 32'h1a712c23;        \
    mem_reg[315] = 32'h01400313;        \
    mem_reg[316] = 32'h00000413;        \
    mem_reg[317] = 32'h408303b3;        \
    mem_reg[318] = 32'h1a712e23;        \
    mem_reg[319] = 32'h00000413;        \
    mem_reg[320] = 32'h406403b3;        \
    mem_reg[321] = 32'h1c712023;        \
    mem_reg[322] = 32'h01900413;        \
    mem_reg[323] = 32'h408303b3;        \
    mem_reg[324] = 32'h1c712223;        \
    mem_reg[325] = 32'hfe700413;        \
    mem_reg[326] = 32'h408303b3;        \
    mem_reg[327] = 32'h1c712423;        \
    mem_reg[328] = 32'h00100313;        \
    mem_reg[329] = 32'h00000413;        \
    mem_reg[330] = 32'h00630463;        \
    mem_reg[331] = 32'h1c812623;        \
    mem_reg[332] = 32'h1c612623;        \
    mem_reg[333] = 32'h14640863;        \
    mem_reg[334] = 32'h1c612823;        \
    mem_reg[335] = 32'h00100313;        \
    mem_reg[336] = 32'h00000413;        \
    mem_reg[337] = 32'h00831463;        \
    mem_reg[338] = 32'h1c812a23;        \
    mem_reg[339] = 32'h1c612a23;        \
    mem_reg[340] = 32'h12631a63;        \
    mem_reg[341] = 32'h1c612c23;        \
    mem_reg[342] = 32'h00600313;        \
    mem_reg[343] = 32'h00700393;        \
    mem_reg[344] = 32'h00800413;        \
    mem_reg[345] = 32'h12634063;        \
    mem_reg[346] = 32'h00734463;        \
    mem_reg[347] = 32'h118001ef;        \
    mem_reg[348] = 32'h10744a63;        \
    mem_reg[349] = 32'h1c612e23;        \
    mem_reg[350] = 32'hff700493;        \
    mem_reg[351] = 32'hff600513;        \
    mem_reg[352] = 32'hff500593;        \
    mem_reg[353] = 32'h1094c063;        \
    mem_reg[354] = 32'h00954463;        \
    mem_reg[355] = 32'h0f8001ef;        \
    mem_reg[356] = 32'h0eb54a63;        \
    mem_reg[357] = 32'h00654463;        \
    mem_reg[358] = 32'h0ec001ef;        \
    mem_reg[359] = 32'h1e612023;        \
    mem_reg[360] = 32'h00600313;        \
    mem_reg[361] = 32'h00700393;        \
    mem_reg[362] = 32'h00800413;        \
    mem_reg[363] = 32'h00635463;        \
    mem_reg[364] = 32'h0d4001ef;        \
    mem_reg[365] = 32'h0063d463;        \
    mem_reg[366] = 32'h0cc001ef;        \
    mem_reg[367] = 32'h0c735463;        \
    mem_reg[368] = 32'h1e612223;        \
    mem_reg[369] = 32'hff700493;        \
    mem_reg[370] = 32'hff600513;        \
    mem_reg[371] = 32'hff500593;        \
    mem_reg[372] = 32'h0094d463;        \
    mem_reg[373] = 32'h0b0001ef;        \
    mem_reg[374] = 32'h00a4d463;        \
    mem_reg[375] = 32'h0a8001ef;        \
    mem_reg[376] = 32'h0aa5d263;        \
    mem_reg[377] = 32'h00935463;        \
    mem_reg[378] = 32'h09c001ef;        \
    mem_reg[379] = 32'h1e612423;        \
    mem_reg[380] = 32'h00600313;        \
    mem_reg[381] = 32'h00700393;        \
    mem_reg[382] = 32'h00800413;        \
    mem_reg[383] = 32'h08636463;        \
    mem_reg[384] = 32'h00736463;        \
    mem_reg[385] = 32'h080001ef;        \
    mem_reg[386] = 32'h06746e63;        \
    mem_reg[387] = 32'h1e612623;        \
    mem_reg[388] = 32'hff700493;        \
    mem_reg[389] = 32'hff600513;        \
    mem_reg[390] = 32'hff500593;        \
    mem_reg[391] = 32'h0694e463;        \
    mem_reg[392] = 32'h00956463;        \
    mem_reg[393] = 32'h060001ef;        \
    mem_reg[394] = 32'h04b56e63;        \
    mem_reg[395] = 32'h04656c63;        \
    mem_reg[396] = 32'h1e612823;        \
    mem_reg[397] = 32'h00600313;        \
    mem_reg[398] = 32'h00700393;        \
    mem_reg[399] = 32'h00800413;        \
    mem_reg[400] = 32'h00637463;        \
    mem_reg[401] = 32'h040001ef;        \
    mem_reg[402] = 32'h0063f463;        \
    mem_reg[403] = 32'h038001ef;        \
    mem_reg[404] = 32'h02737a63;        \
    mem_reg[405] = 32'h1e612a23;        \
    mem_reg[406] = 32'hff700493;        \
    mem_reg[407] = 32'hff600513;        \
    mem_reg[408] = 32'hff500593;        \
    mem_reg[409] = 32'h0094f463;        \
    mem_reg[410] = 32'h01c001ef;        \
    mem_reg[411] = 32'h00a4f463;        \
    mem_reg[412] = 32'h014001ef;        \
    mem_reg[413] = 32'h00a5f863;        \
    mem_reg[414] = 32'h00937663;        \
    mem_reg[415] = 32'h1e612c23;        \
    mem_reg[416] = 32'h000001ef;        \
    mem_reg[417] = 32'h000001ef;

`endif // RISCV_SINGLE_ALL_INSTR_MEM_MAP_SVH