`ifndef ALU_H
`define ALU_H

localparam alu_op_add = 2'b00;
localparam alu_op_sub = 2'b01;
localparam alu_op_and = 2'b10;
localparam alu_op_or  = 2'b11;

`endif // ALU_H