`ifndef MEM_MAP_SVH
`define MEM_MAP_SVH

`define SEC_DATA_W  508

`endif // MEM_MAP_SVH